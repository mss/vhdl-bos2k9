-----------------------------------------------------------------------
-- Copyright (c) 2009 Malte S. Stretz <http://msquadrat.de> 
--
-- TODO: description

-----------------------------------------------------------------------
-- This entity is part of the following library:
-- pragma library fhw_sd
library fhw_sd;
use fhw_sd.sd_globals.all;

library fhw_spi;
use fhw_spi.spi_master;

library fhw_tools;
use fhw_tools.types.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sd_manager_e is
  port(
    clock : in std_logic;
    reset : in std_logic;
    
    address : in std_logic_block_address_t;
    start   : in std_logic;
    
    ready : out std_logic;
    busy  : out std_logic;
    error : out std_logic;
    
    command  : out std_logic_cmd_t;
    argument : out std_logic_arg_t;
    --trigger  : out std_logic;
    shifting : in  std_logic;
    response : in  std_logic_rsp_t);
end sd_manager_e;

-----------------------------------------------------------------------

architecture rtl of sd_manager_e is
  
  type state_t is (
    rset_state_c,
    strt_state_c,
    init_state_c,
    bsiz_state_c,
    read_state_c,
    send_state_c,
    shft_state_c,
    vrfy_state_c,
    idle_state_c);
  signal curr_state_s : state_t;
  signal prev_state_s : state_t;
  signal next_state_s : state_t;
  
  signal error_s : std_logic;

begin
  
  sequence : process(clock, reset)
  begin
    if reset = '1' then
      curr_state_s <= rset_state_c;
    elsif rising_edge(clock) then
      case curr_state_s is
        when rset_state_c => curr_state_s <= strt_state_c;
        when strt_state_c => curr_state_s <= send_state_c;
        when init_state_c => curr_state_s <= send_state_c;
        when bsiz_state_c => curr_state_s <= send_state_c;
        when read_state_c => curr_state_s <= send_state_c;
        when send_state_c => curr_state_s <= shft_state_c;
        when shft_state_c => curr_state_s <= next_state_s;
        when vrfy_state_c => curr_state_s <= next_state_s;
        when idle_state_c => curr_state_s <= next_state_s;
      end case;
    end if;
  end process;
  
  output : process(clock, reset)
    variable address_v : std_logic_arg_t;
  begin
    if rising_edge(clock) then
      prev_state_s <= curr_state_s;
      case curr_state_s is
        when rset_state_c =>
          command  <= cmd_do_reset_c;
          argument <= arg_do_reset_c;
        when strt_state_c =>
          command  <= cmd_do_start_c;
          argument <= arg_do_start_c;
        when init_state_c =>
          command  <= cmd_go_idle_state_c;
          argument <= arg_go_idle_state_c;
        when bsiz_state_c =>
          command  <= cmd_set_blocklen_c;
          argument <= arg_set_blocklen_c;
        when read_state_c =>
          command  <= cmd_read_single_block_c;
          argument <= address & pad_read_single_block_c;
        when others =>
          prev_state_s <= prev_state_s;
      end case;
    end if;
  end process;
  
  -- verify : process(clock, reset, curr_state_s)
  -- begin
    -- if reset = '1' then
      -- error_s <= '0';
    -- elsif rising_edge(clock) then
      -- case curr_state_s is
        -- when shft_state_c =>
          -- if shifting = '0' then
            -- next_state_s <= vrfy_state_c;
          -- end if;
        -- when vrfy_state_c then
          -- if response = "00000000" then
            -- error_s <= '0';
          -- end if;
      -- end case;
    -- end if;
  -- end;
  
  
  
  -- sequence : process(clock, reset, curr_s, next_s)
  -- begin
    -- if error = '1' then
      -- next_s <= rset_state_c;
    -- else
      -- if curr_s = 
    -- end if;
    
    -- case curr_s is
      -- when rset_state_c =>
        -- next_s <= 
    -- end case;
  -- end;
  
  -- output : process(clock, reset, curr_s, next_s)
  -- begin
    
  -- end;
  
  -- transition : process(clock, reset, curr_s, next_s)
  -- begin
    -- if reset = '1' then
      -- curr_s <= reset_state_c;
    -- elsif rising_edge(clock) then
      -- curr_s <= next_s;
    -- end if;
  -- end;
  
end rtl;
